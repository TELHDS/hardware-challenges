// Reference implementation for 8-bit Ripple Carry Adder
// This is a basic implementation for comparison purposes
// Miners should strive to optimize beyond this baseline

module adder_8bit (
    input [7:0] a,
    input [7:0] b, 
    input cin,
    output [7:0] sum,
    output cout
);

    // Internal carry signals
    wire [7:0] carry;
    
    // Full adder for bit 0
    full_adder fa0 (
        .a(a[0]),
        .b(b[0]),
        .cin(cin),
        .sum(sum[0]),
        .cout(carry[0])
    );
    
    // Full adders for bits 1-6
    genvar i;
    generate
        for (i = 1; i < 7; i = i + 1) begin : fa_gen
            full_adder fa (
                .a(a[i]),
                .b(b[i]),
                .cin(carry[i-1]),
                .sum(sum[i]),
                .cout(carry[i])
            );
        end
    endgenerate
    
    // Full adder for bit 7 (MSB)
    full_adder fa7 (
        .a(a[7]),
        .b(b[7]),
        .cin(carry[6]),
        .sum(sum[7]),
        .cout(cout)
    );

endmodule

// Basic full adder module
module full_adder (
    input a,
    input b,
    input cin,
    output sum,
    output cout
);

    // Sum: XOR of all inputs
    assign sum = a ^ b ^ cin;
    
    // Carry: majority function
    assign cout = (a & b) | (cin & (a ^ b));

endmodule
